----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Mike Field <hamster@sanp.net.nz> 
-- 
-- Description: Register settings for the OV7670 Caamera (partially from OV7670.c
--              in the Linux Kernel
------------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ov7670_registers is
    Port ( clk      : in  STD_LOGIC;
           resend   : in  STD_LOGIC;
           advance  : in  STD_LOGIC;
           command  : out  std_logic_vector(15 downto 0);
           finished : out  STD_LOGIC);
end ov7670_registers;

architecture Behavioral of ov7670_registers is
	signal sreg   : std_logic_vector(15 downto 0);
	signal address : std_logic_vector(7 downto 0) := (others => '0');
begin
	command <= sreg;
	with sreg select finished  <= '1' when x"FFFF", '0' when others;
	
	process(clk)
	begin
		if rising_edge(clk) then
			if resend = '1' then 
				address <= (others => '0');
			elsif advance = '1' then
				address <= std_logic_vector(unsigned(address)+1);
			end if;

			case address is
			-- QCIF
				when x"00" => sreg <= x"1280"; -- COM7   Reset
				when x"01" => sreg <= x"1280"; -- COM7   Reset

				when x"02" => sreg <= x"1101"; -- CLKRC
				when x"03" => sreg <= x"1200"; -- COM7
				when x"04" => sreg <= x"0C0C"; -- COM3
				when x"05" => sreg <= x"3E11"; -- COM14
				when x"06" => sreg <= x"703A"; -- SCALING_XSC
				when x"07" => sreg <= x"7135"; -- SCALING_YSC
				when x"08" => sreg <= x"7211"; -- SCALING_DCWCTR
				when x"09" => sreg <= x"73F1"; -- SCALING_PCLK_DIV
				when x"0A" => sreg <= x"A252"; -- SCALING_PCLK_DELAY

-- Attempt to simplify
--				when x"00" => sreg <= x"1280"; -- COM7   Reset
--				when x"01" => sreg <= x"1280"; -- COM7   Reset
--				when x"02" => sreg <= x"1100"; -- CLKRC  Prescaler - Fin/(1+1)
--				when x"03" => sreg <= x"1208"; -- COM7 	 Set format to QCIF 
--				when x"04" => sreg <= x"0C04"; -- COM3  Lots of stuff, enable scaling, all others off
--				when x"05" => sreg <= x"3E19"; -- COM14  PCLK scaling = 0
-- Old Configuration
--				when x"00" => sreg <= x"1280"; -- COM7   Reset
--				when x"01" => sreg <= x"1280"; -- COM7   Reset
--				when x"02" => sreg <= x"1200"; -- COM7   Size & YUV output
--				when x"03" => sreg <= x"1100"; -- CLKRC  Prescaler - Fin/(1+1)
--				when x"04" => sreg <= x"0C00"; -- COM3   Lots of stuff, enable scaling, all others off
--				when x"05" => sreg <= x"3E00"; -- COM14  PCLK scaling off
--				
--				when x"06" => sreg <= x"8C00"; -- RGB444 Set RGB format
--				when x"07" => sreg <= x"0400"; -- COM1   no CCIR601
--				when x"08" => sreg <= x"40C0"; -- COM15  Full 0-255 output
--				when x"09" => sreg <= x"3a00"; -- TSLB   Set UV ordering,  do not auto-reset window
--				when x"0A" => sreg <= x"1438"; -- COM9  - AGC Celling
--				when x"0B" => sreg <= x"4fb3"; -- MTX1  - colour conversion matrix
--				when x"0C" => sreg <= x"50b3"; -- MTX2  - colour conversion matrix
--				when x"0D" => sreg <= x"5100"; -- MTX3  - colour conversion matrix
--				when x"0E" => sreg <= x"523d"; -- MTX4  - colour conversion matrix
--				when x"0F" => sreg <= x"53a7"; -- MTX5  - colour conversion matrix
--				when x"10" => sreg <= x"54e4"; -- MTX6  - colour conversion matrix
--				when x"11" => sreg <= x"589e"; -- MTXS  - Matrix sign and auto contrast
--				when x"12" => sreg <= x"3dc0"; -- COM13 - Turn on GAMMA and UV Auto adjust
--				when x"13" => sreg <= x"1100"; -- CLKRC  Prescaler - Fin/(1+1)
--				
--				when x"14" => sreg <= x"1711"; -- HSTART HREF start (high 8 bits)
--				when x"15" => sreg <= x"1861"; -- HSTOP  HREF stop (high 8 bits)
--				when x"16" => sreg <= x"32A4"; -- HREF   Edge offset and low 3 bits of HSTART and HSTOP
--				
--				when x"17" => sreg <= x"1903"; -- VSTART VSYNC start (high 8 bits)
--				when x"18" => sreg <= x"1A7b"; -- VSTOP  VSYNC stop (high 8 bits) 
--				when x"19" => sreg <= x"030a"; -- VREF   VSYNC low two bits
--				
--				when x"10" => sreg <= x"703a"; -- SCALING_XSC
--				when x"11" => sreg <= x"7135"; -- SCALING_YSC
--				when x"12" => sreg <= x"7200"; -- SCALING_DCWCTR  -- zzz was 11 
--				when x"13" => sreg <= x"7300"; -- SCALING_PCLK_DIV
--				when x"14" => sreg <= x"a200"; -- SCALING_PCLK_DELAY  must match COM14
--          	when x"15" => sreg <= x"1500"; -- COM10 Use HREF not hSYNC
--				
--				when x"1D" => sreg <= x"B104"; -- ABLC1 - Turn on auto black level
--				when x"1F" => sreg <= x"138F"; -- COM8  - AGC, White balance
--				when x"21" => sreg <= x"FFFF"; -- spare
--				when x"22" => sreg <= x"FFFF"; -- spare
--				when x"23" => sreg <= x"0000"; -- spare
--				when x"24" => sreg <= x"0000"; -- spare
--				when x"25" => sreg <= x"138F"; -- COM8 - AGC, White balance
--				when x"26" => sreg <= x"0000"; -- spare
--				when x"27" => sreg <= x"1000"; -- AECH Exposure
--				when x"28" => sreg <= x"0D40"; -- COMM4 - Window Size
--				when x"29" => sreg <= x"0000"; -- spare
--				when x"2a" => sreg <= x"a505"; -- AECGMAX banding filter step
--				when x"2b" => sreg <= x"2495"; -- AEW AGC Stable upper limite
--				when x"2c" => sreg <= x"2533"; -- AEB AGC Stable lower limi
--				when x"2d" => sreg <= x"26e3"; -- VPT AGC fast mode limits
--				when x"2e" => sreg <= x"9f78"; -- HRL High reference level
--				when x"2f" => sreg <= x"A068"; -- LRL low reference level
--				when x"30" => sreg <= x"a103"; -- DSPC3 DSP control
--				when x"31" => sreg <= x"A6d8"; -- LPH Lower Prob High
--				when x"32" => sreg <= x"A7d8"; -- UPL Upper Prob Low
--				when x"33" => sreg <= x"A8f0"; -- TPL Total Prob Low
--				when x"34" => sreg <= x"A990"; -- TPH Total Prob High
--				when x"35" => sreg <= x"AA94"; -- NALG AEC Algo select
--				when x"36" => sreg <= x"13E5"; -- COM8 AGC Settings
				when others => sreg <= x"ffff";
			end case;
		end if;
	end process;
end Behavioral;

